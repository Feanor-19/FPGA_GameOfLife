bind vga asrt_vga asrt_vga_inst (.*);
