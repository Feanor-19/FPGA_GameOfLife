bind vga            asrt_vga            asrt_vga_inst               (.*);
bind NFI_controller asrt_NFI_controller asrt_NFI_controller_inst    (.*);
bind FCL_controller asrt_FCL_controller asrt_FCL_controller_inst    (.*);
