`timescale 1ns/1ps

package defs;

typedef enum logic { FIELD_A, FIELD_B } cur_field_t;
    
endpackage
