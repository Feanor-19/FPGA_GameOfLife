`timescale 1ns/1ps

module tb_get_nbrs_address;

localparam FIELD_W = 4;
localparam FIELD_H = 3;

