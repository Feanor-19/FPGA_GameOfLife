`timescale 1ns/1ps

package defs;

typedef enum logic { 
    FIELD_A, 
    FIELD_B 
} field_t;

typedef enum logic { 
    NO_REQ, 
    CFG_1
} load_cfg_req_t;     

endpackage
